Diente_de_Sierra_inst : Diente_de_Sierra PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
